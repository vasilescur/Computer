`include "../components/mux.v"
`include "../components/mux_thicc.v"
`include "../components/demux.v"
`include "../components/demux_thicc.v"

`include "../components/comparator.v"
`include "../components/adder.v"

`include "../components/ram.v"
`include "../components/rom.v"
`include "../components/register.v"

`include "../components/tty.v"

module computer ();
